module Fetch (
     
);
    
endmodule