module ALU #(
    parameters
) (
    input 
    output
);
    
endmodule