module Immediate_Generator #(
    parameter data_width = 32
) (
    input clk,
    input [data_width-1:0] address
);


    
endmodule